module top (
         input  BTN0
        ,output LED0_G
    ) ;

    assign LED0_G = BTN0 ;

endmodule
